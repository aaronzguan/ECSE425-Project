--********************************************************************
-- ECSE 425, Group 6
-- Kristin Lee (260509976)
-- Date: March 13, 2017

-- Description: ALU_control.vhd

--********************************************************************

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ALU_control is
  port(
      );
end ALU_control;

architecture behaviour of ALU_control is

  begin
  
end behaviour;
